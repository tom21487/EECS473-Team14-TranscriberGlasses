//Copyright (C)2014-2020 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.6.02Beta
//Part Number: GW1NSR-LV4CQN48PC6/I5
//Created Time: Mon Nov 27 14:41:53 2023

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [63:0] dout;
input clk;
input oce;
input ce;
input reset;
input [5:0] ad;

wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO(dout[31:0]),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,gw_gnd,gw_gnd,ad[5:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 32;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0303663C1E16467F1E16467F6666361F0303663C3E66663F33331E0C00000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h6363361C7B6F67637F7F77630606060F1E366667303030780C0C0C1E3F333333;
defparam prom_inst_0.INIT_RAM_02 = 256'h6B63636333333333333333330C0C2D3F0E07331E3E66663F3333331E3E66663F;
defparam prom_inst_0.INIT_RAM_03 = 256'h33363C381C30331E1C30331E0C0C0E0C7B73633E1831637F1E3333331C366363;
defparam prom_inst_0.INIT_RAM_04 = 256'h1830331E00000000000000003E33331E1E33331E1830333F1F03061C301F033F;
defparam prom_inst_0.INIT_RAM_05 = 256'h000C0C003333331E181818183F00000000000000180C06030C183060183C3C18;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000030606;

pROM prom_inst_1 (
    .DO(dout[63:32]),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,gw_gnd,gw_gnd,ad[5:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 32;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h007C6673000F0616007F4616001F3666003C6603003F66660033333F00000000;
defparam prom_inst_1.INIT_RAM_01 = 256'h001C3663006363730063636B007F664600676636001E3333001E0C0C00333333;
defparam prom_inst_1.INIT_RAM_02 = 256'h0063777F000C1E33003F3333001E0C0C001E33380067663600381E3B000F0606;
defparam prom_inst_1.INIT_RAM_03 = 256'h0078307F001E3330003F3306003F0C0C003E676F007F664C001E0C0C0063361C;
defparam prom_inst_1.INIT_RAM_04 = 256'h000C000C060C0C00000C0C00000E1830001E3333000C0C0C001E3333001E3330;
defparam prom_inst_1.INIT_RAM_05 = 256'h000C0C000000001E001818180000000000FF0000004060300001030600180018;
defparam prom_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //Gowin_pROM
