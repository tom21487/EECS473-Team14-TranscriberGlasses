// TODO: port over the fonts here: https://github.com/dhepper/font8x8
`define FONT_BITMAPS \
wire [64*64-1:0] a_bitmap = { \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000000000000000000000000000000000000000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111110000000000011111111111111111111111111111100000000000111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111  \
}; \
wire [64*64-1:0] b_bitmap = { \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111100000000000000000000000000000000000000000000000001111111111, \
    64'b 1111100000000000000000000000000000000000000000000000000011111111, \
    64'b 1111100000000000000000000000000000000000000000000000000011111111, \
    64'b 1111100000000000000000000000000000000000000000000000000011111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000011111111, \
    64'b 1111100000000000000000000000000000000000000000000000000011111111, \
    64'b 1111100000000000000000000000000000000000000000000001111111111111, \
    64'b 1111100000000000000000000000000000000000000000111111111111111111, \
    64'b 1111100000000000000000000000000000000111111111111111111111111111, \
    64'b 1111100000000000000000000000000000011111111111111111111111111111, \
    64'b 1111100000000000000000000000000000000111111111111111111111111111, \
    64'b 1111100000000000000000000000000000000000000000111111111111111111, \
    64'b 1111100000000000000000000000000000000000000000000011111111111111, \
    64'b 1111100000000000000000000000000000000000000000000011111111111111, \
    64'b 1111100000000000000000000000000000000000000000000001111111111111, \
    64'b 1111100000000000000000000000000000000000000000000000000011111111, \
    64'b 1111100000000000011111111111111111111111111111000000000000111111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000001111111, \
    64'b 1111100000000000000000000000000000000000000000000000000011111111, \
    64'b 1111100000000000000000000000000000000000000000000000111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111  \
}; \
wire [64*64-1:0] c_bitmap = { \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111110000000000011111, \
    64'b 1111100000000000011111111111111111111111111111110000000000011111, \
    64'b 1111100000000000011111111111111111111111111111110000000000011111, \
    64'b 1111100000000000011111111111111111111111111111110000000000011111, \
    64'b 1111100000000000011111111111111111111111111111110000000000011111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111000000000001111, \
    64'b 1111100000000000011111111111111111111111111111111000000000001111, \
    64'b 1111100000000000011111111111111111111111111111111000000000001111, \
    64'b 1111100000000000011111111111111111111111111111111000000000001111, \
    64'b 1111100000000000011111111111111111111111111111111000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111  \
}; \
wire [64*64-1:0] d_bitmap = { \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \ 
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111100000000000000000000000000000000000000000000000011111111111, \
    64'b 1111100000000000000000000000000000000000000000000000000001111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000011111111111111111111111111111100000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000001111111, \
    64'b 1111100000000000000000000000000000000000000000000000000011111111, \
    64'b 1111100000000000000000000000000000000000000000000000001111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111  \
}; \
wire [64*64-1:0] e_bitmap = { \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000000000000000000000000000000000000000000000011111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000011111111111111111111111111111111111111111111111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111100000000000000000000000000000000000000000000000000000001111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111, \
    64'b 1111111111111111111111111111111111111111111111111111111111111111  \
};
